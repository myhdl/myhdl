module const_1(q, clk);

   input clk;
   output q;

   wire q = 1;

endmodule // inc
